/*Mux
---------------------------------------------------------
| S | A | B | Y |				   
|---------------|				      S
| 0   0   0   0	|				      |
|---------------|				 _____|____
| 0   0   1   1 |				|	  	   \
|---------------|				|  Mux	   |
| 0   1   0   0 |				|	  	   |
|---------------|		   A----|	       |
| 0   1   1   1 |				|	  	   |----Y
|_______________|				|	       |
|_______________|				|	  	   |
| 1   0   0   0 |				|	       |
|---------------|		   B----|	  	   |
| 1   0   1   0 |				|	       |
|---------------|				|_________/
| 1   1   0   1 |
|---------------|
| 1   1   1   1 |
---------------------------------------------------------
*/
module Mux2ver (
	input wire Select,	       // the switching signal
    input wire A_in,	       // input line
	input wire B_in,	       // input line

    output Y			   // output line	
);

assign Y = (Select) ? A_in : B_in;
endmodule
